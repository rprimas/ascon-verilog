logic [127:0] tb_key = 128'h0F0E0D0C0B0A09080706050403020100;
logic [127:0] tb_nonce = 128'h0F0E0D0C0B0A09080706050403020100;
logic [127:0] tb_tag = 128'h732ED5035140D9B19B2520E2E36C3A86;
logic [31:0] tb_ad = 32'h03020100;
logic [31:0] tb_msg = 32'h03020100;
logic [31:0] tb_ct = 32'h96D9534A;
logic [255:0] tb_hash = 256'hEE2767DF377184FDD7B2E14F30D8EC547087F859F29E8BD05C328A9BEDC7E4D7;
